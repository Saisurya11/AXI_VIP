// Code your testbench here
// or browse Examples
`include "axi_top.sv"